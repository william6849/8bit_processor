module PC_add(a,b,out);
	input [4:0]a,b;
	output [4:0]out;

	assign out=a+b;

endmodule